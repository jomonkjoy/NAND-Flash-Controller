module nand_flash_controller #(
) (
);

endmodule
